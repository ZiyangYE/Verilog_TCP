function logic [31:0] compute_crc_16(input [31:0] crc_reg, input [127:0] data_in);
    logic [31:0] crc_out;

    crc_out[31] = crc_reg[31] ^ crc_reg[30] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[26] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[21] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[4] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[1] ^ data_in[14] ^ data_in[13] ^ data_in[11] ^ data_in[23] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[39] ^ data_in[37] ^ data_in[34] ^ data_in[43] ^ data_in[42] ^ data_in[40] ^ data_in[55] ^ data_in[53] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[61] ^ data_in[59] ^ data_in[58] ^ data_in[56] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[79] ^ data_in[78] ^ data_in[72] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[80] ^ data_in[89] ^ data_in[88] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[98] ^ data_in[96] ^ data_in[111] ^ data_in[109] ^ data_in[105] ^ data_in[104] ^ data_in[118] ^ data_in[117] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[124] ^ data_in[122] ^ data_in[121] ^ data_in[120];
    crc_out[30] = crc_reg[27] ^ crc_reg[26] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[17] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[7] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[7] ^ data_in[6] ^ data_in[1] ^ data_in[0] ^ data_in[14] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[23] ^ data_in[22] ^ data_in[31] ^ data_in[28] ^ data_in[27] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[34] ^ data_in[33] ^ data_in[43] ^ data_in[41] ^ data_in[40] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[50] ^ data_in[63] ^ data_in[61] ^ data_in[60] ^ data_in[59] ^ data_in[57] ^ data_in[56] ^ data_in[71] ^ data_in[70] ^ data_in[66] ^ data_in[79] ^ data_in[77] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[81] ^ data_in[80] ^ data_in[95] ^ data_in[89] ^ data_in[99] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[105] ^ data_in[119] ^ data_in[118] ^ data_in[116] ^ data_in[115] ^ data_in[127] ^ data_in[124] ^ data_in[123] ^ data_in[122];
    crc_out[29] = crc_reg[31] ^ crc_reg[30] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[25] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[17] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[1] ^ data_in[0] ^ data_in[15] ^ data_in[14] ^ data_in[10] ^ data_in[9] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[31] ^ data_in[29] ^ data_in[25] ^ data_in[24] ^ data_in[39] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[43] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[48] ^ data_in[62] ^ data_in[61] ^ data_in[60] ^ data_in[71] ^ data_in[68] ^ data_in[67] ^ data_in[65] ^ data_in[79] ^ data_in[76] ^ data_in[72] ^ data_in[87] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[95] ^ data_in[94] ^ data_in[89] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[97] ^ data_in[108] ^ data_in[107] ^ data_in[105] ^ data_in[113] ^ data_in[112] ^ data_in[126] ^ data_in[124] ^ data_in[123] ^ data_in[120];
    crc_out[28] = crc_reg[30] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[24] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[16] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[0] ^ data_in[15] ^ data_in[14] ^ data_in[13] ^ data_in[9] ^ data_in[8] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[30] ^ data_in[28] ^ data_in[24] ^ data_in[39] ^ data_in[38] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[47] ^ data_in[42] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[63] ^ data_in[61] ^ data_in[60] ^ data_in[59] ^ data_in[70] ^ data_in[67] ^ data_in[66] ^ data_in[64] ^ data_in[78] ^ data_in[75] ^ data_in[87] ^ data_in[86] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[94] ^ data_in[93] ^ data_in[88] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[96] ^ data_in[107] ^ data_in[106] ^ data_in[104] ^ data_in[112] ^ data_in[127] ^ data_in[125] ^ data_in[123] ^ data_in[122];
    crc_out[27] = crc_reg[30] ^ crc_reg[27] ^ crc_reg[24] ^ crc_reg[21] ^ crc_reg[18] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[0] ^ data_in[7] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[1] ^ data_in[15] ^ data_in[12] ^ data_in[11] ^ data_in[8] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[31] ^ data_in[30] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[38] ^ data_in[33] ^ data_in[32] ^ data_in[47] ^ data_in[46] ^ data_in[43] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[55] ^ data_in[53] ^ data_in[62] ^ data_in[61] ^ data_in[60] ^ data_in[56] ^ data_in[70] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[78] ^ data_in[77] ^ data_in[74] ^ data_in[72] ^ data_in[84] ^ data_in[83] ^ data_in[81] ^ data_in[93] ^ data_in[92] ^ data_in[89] ^ data_in[88] ^ data_in[102] ^ data_in[99] ^ data_in[96] ^ data_in[109] ^ data_in[106] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[120];
    crc_out[26] = crc_reg[30] ^ crc_reg[28] ^ crc_reg[24] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ^ data_in[13] ^ data_in[10] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[31] ^ data_in[27] ^ data_in[26] ^ data_in[34] ^ data_in[32] ^ data_in[47] ^ data_in[46] ^ data_in[45] ^ data_in[43] ^ data_in[41] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[60] ^ data_in[58] ^ data_in[56] ^ data_in[71] ^ data_in[70] ^ data_in[68] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[73] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[92] ^ data_in[91] ^ data_in[89] ^ data_in[102] ^ data_in[100] ^ data_in[96] ^ data_in[109] ^ data_in[108] ^ data_in[104] ^ data_in[119] ^ data_in[116] ^ data_in[115] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[122] ^ data_in[121] ^ data_in[120];
    crc_out[25] = crc_reg[29] ^ crc_reg[27] ^ crc_reg[23] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ^ data_in[15] ^ data_in[12] ^ data_in[9] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[30] ^ data_in[26] ^ data_in[25] ^ data_in[33] ^ data_in[47] ^ data_in[46] ^ data_in[45] ^ data_in[44] ^ data_in[42] ^ data_in[40] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[49] ^ data_in[48] ^ data_in[63] ^ data_in[59] ^ data_in[57] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[67] ^ data_in[65] ^ data_in[64] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[91] ^ data_in[90] ^ data_in[88] ^ data_in[101] ^ data_in[99] ^ data_in[111] ^ data_in[108] ^ data_in[107] ^ data_in[119] ^ data_in[118] ^ data_in[115] ^ data_in[114] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[121] ^ data_in[120];
    crc_out[24] = crc_reg[30] ^ crc_reg[29] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[11] ^ crc_reg[8] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[1] ^ data_in[7] ^ data_in[5] ^ data_in[4] ^ data_in[2] ^ data_in[0] ^ data_in[15] ^ data_in[13] ^ data_in[8] ^ data_in[23] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[31] ^ data_in[30] ^ data_in[27] ^ data_in[26] ^ data_in[39] ^ data_in[37] ^ data_in[34] ^ data_in[32] ^ data_in[46] ^ data_in[45] ^ data_in[44] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[49] ^ data_in[63] ^ data_in[62] ^ data_in[61] ^ data_in[59] ^ data_in[67] ^ data_in[66] ^ data_in[64] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[72] ^ data_in[87] ^ data_in[80] ^ data_in[90] ^ data_in[88] ^ data_in[102] ^ data_in[101] ^ data_in[96] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[115] ^ data_in[112] ^ data_in[125] ^ data_in[123] ^ data_in[121];
    crc_out[23] = crc_reg[30] ^ crc_reg[26] ^ crc_reg[24] ^ crc_reg[22] ^ crc_reg[20] ^ crc_reg[18] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[11] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[1] ^ data_in[7] ^ data_in[6] ^ data_in[4] ^ data_in[3] ^ data_in[15] ^ data_in[13] ^ data_in[12] ^ data_in[11] ^ data_in[22] ^ data_in[17] ^ data_in[16] ^ data_in[27] ^ data_in[24] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[34] ^ data_in[33] ^ data_in[47] ^ data_in[45] ^ data_in[44] ^ data_in[42] ^ data_in[41] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[49] ^ data_in[62] ^ data_in[60] ^ data_in[59] ^ data_in[56] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[78] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[87] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[80] ^ data_in[95] ^ data_in[88] ^ data_in[102] ^ data_in[98] ^ data_in[96] ^ data_in[110] ^ data_in[108] ^ data_in[106] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[115] ^ data_in[113] ^ data_in[112] ^ data_in[127] ^ data_in[121];
    crc_out[22] = crc_reg[31] ^ crc_reg[29] ^ crc_reg[25] ^ crc_reg[23] ^ crc_reg[21] ^ crc_reg[19] ^ crc_reg[17] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[3] ^ data_in[2] ^ data_in[14] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[21] ^ data_in[16] ^ data_in[31] ^ data_in[26] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[33] ^ data_in[32] ^ data_in[46] ^ data_in[44] ^ data_in[43] ^ data_in[41] ^ data_in[40] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[48] ^ data_in[61] ^ data_in[59] ^ data_in[58] ^ data_in[71] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[77] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[95] ^ data_in[94] ^ data_in[103] ^ data_in[101] ^ data_in[97] ^ data_in[111] ^ data_in[109] ^ data_in[107] ^ data_in[105] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[120];
    crc_out[21] = crc_reg[31] ^ crc_reg[29] ^ crc_reg[26] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[14] ^ crc_reg[12] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[5] ^ data_in[4] ^ data_in[2] ^ data_in[14] ^ data_in[10] ^ data_in[9] ^ data_in[23] ^ data_in[20] ^ data_in[29] ^ data_in[27] ^ data_in[26] ^ data_in[24] ^ data_in[39] ^ data_in[38] ^ data_in[36] ^ data_in[35] ^ data_in[32] ^ data_in[47] ^ data_in[45] ^ data_in[53] ^ data_in[51] ^ data_in[48] ^ data_in[63] ^ data_in[61] ^ data_in[60] ^ data_in[59] ^ data_in[57] ^ data_in[56] ^ data_in[69] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[78] ^ data_in[76] ^ data_in[74] ^ data_in[73] ^ data_in[87] ^ data_in[84] ^ data_in[81] ^ data_in[94] ^ data_in[93] ^ data_in[89] ^ data_in[88] ^ data_in[103] ^ data_in[101] ^ data_in[98] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[106] ^ data_in[105] ^ data_in[118] ^ data_in[116] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[122] ^ data_in[121] ^ data_in[120];
    crc_out[20] = crc_reg[29] ^ crc_reg[26] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[14] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[7] ^ data_in[6] ^ data_in[4] ^ data_in[3] ^ data_in[14] ^ data_in[11] ^ data_in[9] ^ data_in[8] ^ data_in[23] ^ data_in[22] ^ data_in[19] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[24] ^ data_in[38] ^ data_in[35] ^ data_in[47] ^ data_in[46] ^ data_in[44] ^ data_in[43] ^ data_in[42] ^ data_in[40] ^ data_in[55] ^ data_in[53] ^ data_in[52] ^ data_in[49] ^ data_in[48] ^ data_in[63] ^ data_in[62] ^ data_in[61] ^ data_in[60] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[67] ^ data_in[65] ^ data_in[64] ^ data_in[78] ^ data_in[77] ^ data_in[75] ^ data_in[73] ^ data_in[85] ^ data_in[84] ^ data_in[82] ^ data_in[93] ^ data_in[92] ^ data_in[89] ^ data_in[101] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[111] ^ data_in[110] ^ data_in[108] ^ data_in[107] ^ data_in[118] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[123] ^ data_in[122];
    crc_out[19] = crc_reg[31] ^ crc_reg[30] ^ crc_reg[29] ^ crc_reg[26] ^ crc_reg[25] ^ crc_reg[22] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[14] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[14] ^ data_in[11] ^ data_in[10] ^ data_in[8] ^ data_in[22] ^ data_in[21] ^ data_in[18] ^ data_in[31] ^ data_in[28] ^ data_in[25] ^ data_in[24] ^ data_in[46] ^ data_in[45] ^ data_in[41] ^ data_in[40] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[63] ^ data_in[62] ^ data_in[60] ^ data_in[58] ^ data_in[56] ^ data_in[67] ^ data_in[66] ^ data_in[64] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[74] ^ data_in[86] ^ data_in[85] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[92] ^ data_in[91] ^ data_in[89] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[98] ^ data_in[97] ^ data_in[110] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[118] ^ data_in[115] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[120];
    crc_out[18] = crc_reg[30] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[21] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[13] ^ crc_reg[10] ^ crc_reg[9] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[2] ^ data_in[1] ^ data_in[0] ^ data_in[13] ^ data_in[10] ^ data_in[9] ^ data_in[23] ^ data_in[21] ^ data_in[20] ^ data_in[17] ^ data_in[30] ^ data_in[27] ^ data_in[24] ^ data_in[39] ^ data_in[45] ^ data_in[44] ^ data_in[40] ^ data_in[55] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[62] ^ data_in[61] ^ data_in[59] ^ data_in[57] ^ data_in[71] ^ data_in[66] ^ data_in[65] ^ data_in[79] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[73] ^ data_in[85] ^ data_in[84] ^ data_in[81] ^ data_in[80] ^ data_in[95] ^ data_in[91] ^ data_in[90] ^ data_in[88] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[97] ^ data_in[96] ^ data_in[109] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[119] ^ data_in[117] ^ data_in[114] ^ data_in[113] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124];
    crc_out[17] = crc_reg[31] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[20] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[12] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[1] ^ data_in[0] ^ data_in[15] ^ data_in[12] ^ data_in[9] ^ data_in[8] ^ data_in[22] ^ data_in[20] ^ data_in[19] ^ data_in[16] ^ data_in[29] ^ data_in[26] ^ data_in[39] ^ data_in[38] ^ data_in[44] ^ data_in[43] ^ data_in[55] ^ data_in[54] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[63] ^ data_in[61] ^ data_in[60] ^ data_in[58] ^ data_in[56] ^ data_in[70] ^ data_in[65] ^ data_in[64] ^ data_in[78] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[72] ^ data_in[84] ^ data_in[83] ^ data_in[80] ^ data_in[95] ^ data_in[94] ^ data_in[90] ^ data_in[89] ^ data_in[103] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[96] ^ data_in[111] ^ data_in[108] ^ data_in[105] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[116] ^ data_in[113] ^ data_in[112] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123];
    crc_out[16] = crc_reg[30] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[26] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[19] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[11] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[0] ^ data_in[15] ^ data_in[14] ^ data_in[11] ^ data_in[8] ^ data_in[23] ^ data_in[21] ^ data_in[19] ^ data_in[18] ^ data_in[31] ^ data_in[28] ^ data_in[25] ^ data_in[38] ^ data_in[37] ^ data_in[43] ^ data_in[42] ^ data_in[54] ^ data_in[53] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[63] ^ data_in[62] ^ data_in[60] ^ data_in[59] ^ data_in[57] ^ data_in[71] ^ data_in[69] ^ data_in[64] ^ data_in[79] ^ data_in[77] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[87] ^ data_in[83] ^ data_in[82] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[89] ^ data_in[88] ^ data_in[102] ^ data_in[100] ^ data_in[99] ^ data_in[98] ^ data_in[111] ^ data_in[110] ^ data_in[107] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[115] ^ data_in[112] ^ data_in[127] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[122];
    crc_out[15] = crc_reg[30] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[3] ^ crc_reg[0] ^ data_in[7] ^ data_in[3] ^ data_in[2] ^ data_in[15] ^ data_in[11] ^ data_in[10] ^ data_in[22] ^ data_in[20] ^ data_in[18] ^ data_in[17] ^ data_in[31] ^ data_in[29] ^ data_in[26] ^ data_in[25] ^ data_in[39] ^ data_in[36] ^ data_in[34] ^ data_in[43] ^ data_in[41] ^ data_in[40] ^ data_in[55] ^ data_in[52] ^ data_in[63] ^ data_in[62] ^ data_in[69] ^ data_in[67] ^ data_in[76] ^ data_in[74] ^ data_in[73] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[81] ^ data_in[80] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[89] ^ data_in[102] ^ data_in[100] ^ data_in[99] ^ data_in[97] ^ data_in[96] ^ data_in[111] ^ data_in[110] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[119] ^ data_in[116] ^ data_in[115] ^ data_in[113] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[123] ^ data_in[120];
    crc_out[14] = crc_reg[29] ^ crc_reg[27] ^ crc_reg[26] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[2] ^ data_in[6] ^ data_in[2] ^ data_in[1] ^ data_in[14] ^ data_in[10] ^ data_in[9] ^ data_in[21] ^ data_in[19] ^ data_in[17] ^ data_in[16] ^ data_in[30] ^ data_in[28] ^ data_in[25] ^ data_in[24] ^ data_in[38] ^ data_in[35] ^ data_in[33] ^ data_in[42] ^ data_in[40] ^ data_in[55] ^ data_in[54] ^ data_in[51] ^ data_in[62] ^ data_in[61] ^ data_in[68] ^ data_in[66] ^ data_in[75] ^ data_in[73] ^ data_in[72] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[80] ^ data_in[95] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[88] ^ data_in[101] ^ data_in[99] ^ data_in[98] ^ data_in[96] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[105] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[115] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[122];
    crc_out[13] = crc_reg[31] ^ crc_reg[28] ^ crc_reg[26] ^ crc_reg[25] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[10] ^ crc_reg[9] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[1] ^ data_in[5] ^ data_in[1] ^ data_in[0] ^ data_in[13] ^ data_in[9] ^ data_in[8] ^ data_in[20] ^ data_in[18] ^ data_in[16] ^ data_in[31] ^ data_in[29] ^ data_in[27] ^ data_in[24] ^ data_in[39] ^ data_in[37] ^ data_in[34] ^ data_in[32] ^ data_in[41] ^ data_in[55] ^ data_in[54] ^ data_in[53] ^ data_in[50] ^ data_in[61] ^ data_in[60] ^ data_in[67] ^ data_in[65] ^ data_in[74] ^ data_in[72] ^ data_in[87] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[95] ^ data_in[94] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[103] ^ data_in[100] ^ data_in[98] ^ data_in[97] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[114] ^ data_in[113] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[121];
    crc_out[12] = crc_reg[30] ^ crc_reg[27] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[0] ^ data_in[4] ^ data_in[0] ^ data_in[15] ^ data_in[12] ^ data_in[8] ^ data_in[23] ^ data_in[19] ^ data_in[17] ^ data_in[31] ^ data_in[30] ^ data_in[28] ^ data_in[26] ^ data_in[39] ^ data_in[38] ^ data_in[36] ^ data_in[33] ^ data_in[47] ^ data_in[40] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[49] ^ data_in[60] ^ data_in[59] ^ data_in[66] ^ data_in[64] ^ data_in[73] ^ data_in[87] ^ data_in[86] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[94] ^ data_in[93] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[102] ^ data_in[99] ^ data_in[97] ^ data_in[96] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[107] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[113] ^ data_in[112] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[120];
    crc_out[11] = crc_reg[29] ^ crc_reg[26] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[3] ^ data_in[15] ^ data_in[14] ^ data_in[11] ^ data_in[23] ^ data_in[22] ^ data_in[18] ^ data_in[16] ^ data_in[30] ^ data_in[29] ^ data_in[27] ^ data_in[25] ^ data_in[38] ^ data_in[37] ^ data_in[35] ^ data_in[32] ^ data_in[46] ^ data_in[55] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[48] ^ data_in[59] ^ data_in[58] ^ data_in[65] ^ data_in[79] ^ data_in[72] ^ data_in[86] ^ data_in[85] ^ data_in[81] ^ data_in[80] ^ data_in[95] ^ data_in[93] ^ data_in[92] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[101] ^ data_in[98] ^ data_in[96] ^ data_in[111] ^ data_in[109] ^ data_in[108] ^ data_in[107] ^ data_in[106] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[112] ^ data_in[127] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[122];
    crc_out[10] = crc_reg[31] ^ crc_reg[28] ^ crc_reg[25] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[1] ^ data_in[2] ^ data_in[14] ^ data_in[13] ^ data_in[10] ^ data_in[22] ^ data_in[21] ^ data_in[17] ^ data_in[31] ^ data_in[29] ^ data_in[28] ^ data_in[26] ^ data_in[24] ^ data_in[37] ^ data_in[36] ^ data_in[34] ^ data_in[47] ^ data_in[45] ^ data_in[54] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[63] ^ data_in[58] ^ data_in[57] ^ data_in[64] ^ data_in[78] ^ data_in[87] ^ data_in[85] ^ data_in[84] ^ data_in[80] ^ data_in[95] ^ data_in[94] ^ data_in[92] ^ data_in[91] ^ data_in[89] ^ data_in[88] ^ data_in[103] ^ data_in[100] ^ data_in[97] ^ data_in[111] ^ data_in[110] ^ data_in[108] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[114] ^ data_in[127] ^ data_in[126] ^ data_in[124] ^ data_in[123] ^ data_in[122] ^ data_in[121];
    crc_out[9] = crc_reg[29] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[26] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[8] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ data_in[7] ^ data_in[14] ^ data_in[12] ^ data_in[11] ^ data_in[9] ^ data_in[23] ^ data_in[21] ^ data_in[20] ^ data_in[16] ^ data_in[31] ^ data_in[29] ^ data_in[28] ^ data_in[26] ^ data_in[24] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[46] ^ data_in[44] ^ data_in[43] ^ data_in[42] ^ data_in[40] ^ data_in[55] ^ data_in[51] ^ data_in[48] ^ data_in[62] ^ data_in[61] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[78] ^ data_in[77] ^ data_in[72] ^ data_in[85] ^ data_in[82] ^ data_in[80] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[98] ^ data_in[111] ^ data_in[110] ^ data_in[107] ^ data_in[106] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[112] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123];
    crc_out[8] = crc_reg[31] ^ crc_reg[30] ^ crc_reg[29] ^ crc_reg[27] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[18] ^ crc_reg[16] ^ crc_reg[14] ^ crc_reg[12] ^ crc_reg[10] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[1] ^ data_in[14] ^ data_in[10] ^ data_in[8] ^ data_in[23] ^ data_in[22] ^ data_in[20] ^ data_in[19] ^ data_in[29] ^ data_in[28] ^ data_in[26] ^ data_in[24] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[33] ^ data_in[32] ^ data_in[45] ^ data_in[41] ^ data_in[40] ^ data_in[54] ^ data_in[53] ^ data_in[49] ^ data_in[48] ^ data_in[63] ^ data_in[60] ^ data_in[59] ^ data_in[57] ^ data_in[70] ^ data_in[66] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[90] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[99] ^ data_in[97] ^ data_in[96] ^ data_in[111] ^ data_in[110] ^ data_in[106] ^ data_in[104] ^ data_in[118] ^ data_in[116] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[127] ^ data_in[125] ^ data_in[123] ^ data_in[121] ^ data_in[120];
    crc_out[7] = crc_reg[30] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[26] ^ crc_reg[24] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[17] ^ crc_reg[15] ^ crc_reg[13] ^ crc_reg[11] ^ crc_reg[9] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[2] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[0] ^ data_in[13] ^ data_in[9] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[19] ^ data_in[18] ^ data_in[28] ^ data_in[27] ^ data_in[25] ^ data_in[39] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[32] ^ data_in[47] ^ data_in[44] ^ data_in[40] ^ data_in[55] ^ data_in[53] ^ data_in[52] ^ data_in[48] ^ data_in[63] ^ data_in[62] ^ data_in[59] ^ data_in[58] ^ data_in[56] ^ data_in[69] ^ data_in[65] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[89] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[98] ^ data_in[96] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[105] ^ data_in[119] ^ data_in[117] ^ data_in[115] ^ data_in[113] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[124] ^ data_in[122] ^ data_in[120];
    crc_out[6] = crc_reg[29] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[25] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[16] ^ crc_reg[14] ^ crc_reg[12] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[1] ^ data_in[5] ^ data_in[4] ^ data_in[15] ^ data_in[12] ^ data_in[8] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[18] ^ data_in[17] ^ data_in[27] ^ data_in[26] ^ data_in[24] ^ data_in[38] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[47] ^ data_in[46] ^ data_in[43] ^ data_in[55] ^ data_in[54] ^ data_in[52] ^ data_in[51] ^ data_in[63] ^ data_in[62] ^ data_in[61] ^ data_in[58] ^ data_in[57] ^ data_in[71] ^ data_in[68] ^ data_in[64] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[81] ^ data_in[80] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[88] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[97] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[104] ^ data_in[118] ^ data_in[116] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[123] ^ data_in[121];
    crc_out[5] = crc_reg[30] ^ crc_reg[29] ^ crc_reg[27] ^ crc_reg[23] ^ crc_reg[22] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[10] ^ crc_reg[8] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[1] ^ data_in[7] ^ data_in[4] ^ data_in[3] ^ data_in[1] ^ data_in[13] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[17] ^ data_in[16] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[27] ^ data_in[24] ^ data_in[33] ^ data_in[32] ^ data_in[46] ^ data_in[45] ^ data_in[43] ^ data_in[40] ^ data_in[55] ^ data_in[54] ^ data_in[51] ^ data_in[49] ^ data_in[48] ^ data_in[62] ^ data_in[60] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[69] ^ data_in[68] ^ data_in[78] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[86] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[88] ^ data_in[102] ^ data_in[101] ^ data_in[99] ^ data_in[111] ^ data_in[110] ^ data_in[108] ^ data_in[107] ^ data_in[105] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[114] ^ data_in[112] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[121];
    crc_out[4] = crc_reg[31] ^ crc_reg[29] ^ crc_reg[28] ^ crc_reg[26] ^ crc_reg[22] ^ crc_reg[21] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[9] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[0] ^ data_in[6] ^ data_in[3] ^ data_in[2] ^ data_in[0] ^ data_in[12] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[16] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[26] ^ data_in[39] ^ data_in[32] ^ data_in[47] ^ data_in[45] ^ data_in[44] ^ data_in[42] ^ data_in[55] ^ data_in[54] ^ data_in[53] ^ data_in[50] ^ data_in[48] ^ data_in[63] ^ data_in[61] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[56] ^ data_in[68] ^ data_in[67] ^ data_in[77] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[87] ^ data_in[85] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[103] ^ data_in[101] ^ data_in[100] ^ data_in[98] ^ data_in[110] ^ data_in[109] ^ data_in[107] ^ data_in[106] ^ data_in[104] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[113] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[120];
    crc_out[3] = crc_reg[30] ^ crc_reg[28] ^ crc_reg[27] ^ crc_reg[25] ^ crc_reg[21] ^ crc_reg[20] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[8] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ data_in[5] ^ data_in[2] ^ data_in[1] ^ data_in[15] ^ data_in[11] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[25] ^ data_in[38] ^ data_in[47] ^ data_in[46] ^ data_in[44] ^ data_in[43] ^ data_in[41] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[49] ^ data_in[63] ^ data_in[62] ^ data_in[60] ^ data_in[58] ^ data_in[57] ^ data_in[56] ^ data_in[71] ^ data_in[67] ^ data_in[66] ^ data_in[76] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[84] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[102] ^ data_in[100] ^ data_in[99] ^ data_in[97] ^ data_in[109] ^ data_in[108] ^ data_in[106] ^ data_in[105] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[112] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123];
    crc_out[2] = crc_reg[31] ^ crc_reg[29] ^ crc_reg[27] ^ crc_reg[26] ^ crc_reg[24] ^ crc_reg[20] ^ crc_reg[19] ^ crc_reg[17] ^ crc_reg[16] ^ crc_reg[14] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[7] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[4] ^ data_in[1] ^ data_in[0] ^ data_in[14] ^ data_in[10] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[24] ^ data_in[37] ^ data_in[46] ^ data_in[45] ^ data_in[43] ^ data_in[42] ^ data_in[40] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[48] ^ data_in[62] ^ data_in[61] ^ data_in[59] ^ data_in[57] ^ data_in[56] ^ data_in[71] ^ data_in[70] ^ data_in[66] ^ data_in[65] ^ data_in[75] ^ data_in[73] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[83] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[103] ^ data_in[101] ^ data_in[99] ^ data_in[98] ^ data_in[96] ^ data_in[108] ^ data_in[107] ^ data_in[105] ^ data_in[104] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[127] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[122];
    crc_out[1] = crc_reg[31] ^ crc_reg[30] ^ crc_reg[28] ^ crc_reg[26] ^ crc_reg[25] ^ crc_reg[23] ^ crc_reg[19] ^ crc_reg[18] ^ crc_reg[16] ^ crc_reg[15] ^ crc_reg[13] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[1] ^ data_in[3] ^ data_in[0] ^ data_in[15] ^ data_in[13] ^ data_in[9] ^ data_in[17] ^ data_in[16] ^ data_in[31] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[39] ^ data_in[36] ^ data_in[45] ^ data_in[44] ^ data_in[42] ^ data_in[41] ^ data_in[55] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[63] ^ data_in[61] ^ data_in[60] ^ data_in[58] ^ data_in[56] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[65] ^ data_in[64] ^ data_in[74] ^ data_in[72] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[82] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[103] ^ data_in[102] ^ data_in[100] ^ data_in[98] ^ data_in[97] ^ data_in[111] ^ data_in[107] ^ data_in[106] ^ data_in[104] ^ data_in[119] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[114] ^ data_in[126] ^ data_in[124] ^ data_in[123] ^ data_in[122] ^ data_in[121];
    crc_out[0] = crc_reg[31] ^ crc_reg[30] ^ crc_reg[29] ^ crc_reg[27] ^ crc_reg[25] ^ crc_reg[24] ^ crc_reg[22] ^ crc_reg[18] ^ crc_reg[17] ^ crc_reg[15] ^ crc_reg[14] ^ crc_reg[12] ^ crc_reg[11] ^ crc_reg[10] ^ crc_reg[9] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[2] ^ data_in[15] ^ data_in[14] ^ data_in[12] ^ data_in[8] ^ data_in[16] ^ data_in[31] ^ data_in[30] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[38] ^ data_in[35] ^ data_in[44] ^ data_in[43] ^ data_in[41] ^ data_in[40] ^ data_in[54] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[62] ^ data_in[60] ^ data_in[59] ^ data_in[57] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[64] ^ data_in[79] ^ data_in[73] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[81] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[99] ^ data_in[97] ^ data_in[96] ^ data_in[110] ^ data_in[106] ^ data_in[105] ^ data_in[119] ^ data_in[118] ^ data_in[116] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[125] ^ data_in[123] ^ data_in[122] ^ data_in[121] ^ data_in[120];

    return crc_out;
endfunction

function logic [31:0] compute_crc_1(input [31:0] crc_reg, input [7:0] data_in);
    logic [31:0] crc_out;

    crc_out[31] = crc_reg[7] ^ crc_reg[1] ^ data_in[7] ^ data_in[1];
    crc_out[30] = crc_reg[7] ^ crc_reg[6] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[1] ^ data_in[0];
    crc_out[29] = crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[1] ^ data_in[0];
    crc_out[28] = crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[0];
    crc_out[27] = crc_reg[7] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[1] ^ data_in[7] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[1];
    crc_out[26] = crc_reg[7] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[7] ^ data_in[6] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0];
    crc_out[25] = crc_reg[6] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0];
    crc_out[24] = crc_reg[7] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[2] ^ crc_reg[0] ^ data_in[7] ^ data_in[5] ^ data_in[4] ^ data_in[2] ^ data_in[0];
    crc_out[23] = crc_reg[31] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[3] ^ data_in[7] ^ data_in[6] ^ data_in[4] ^ data_in[3];
    crc_out[22] = crc_reg[30] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[6] ^ data_in[5] ^ data_in[3] ^ data_in[2];
    crc_out[21] = crc_reg[29] ^ crc_reg[7] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[2] ^ data_in[7] ^ data_in[5] ^ data_in[4] ^ data_in[2];
    crc_out[20] = crc_reg[28] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[4] ^ crc_reg[3] ^ data_in[7] ^ data_in[6] ^ data_in[4] ^ data_in[3];
    crc_out[19] = crc_reg[27] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[1] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[3] ^ data_in[2] ^ data_in[1];
    crc_out[18] = crc_reg[26] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[2] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[2] ^ data_in[1] ^ data_in[0];
    crc_out[17] = crc_reg[25] ^ crc_reg[5] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[1] ^ data_in[0];
    crc_out[16] = crc_reg[24] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[0] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[0];
    crc_out[15] = crc_reg[23] ^ crc_reg[7] ^ crc_reg[3] ^ crc_reg[2] ^ data_in[7] ^ data_in[3] ^ data_in[2];
    crc_out[14] = crc_reg[22] ^ crc_reg[6] ^ crc_reg[2] ^ crc_reg[1] ^ data_in[6] ^ data_in[2] ^ data_in[1];
    crc_out[13] = crc_reg[21] ^ crc_reg[5] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[5] ^ data_in[1] ^ data_in[0];
    crc_out[12] = crc_reg[20] ^ crc_reg[4] ^ crc_reg[0] ^ data_in[4] ^ data_in[0];
    crc_out[11] = crc_reg[19] ^ crc_reg[3] ^ data_in[3];
    crc_out[10] = crc_reg[18] ^ crc_reg[2] ^ data_in[2];
    crc_out[9] = crc_reg[17] ^ crc_reg[7] ^ data_in[7];
    crc_out[8] = crc_reg[16] ^ crc_reg[7] ^ crc_reg[6] ^ crc_reg[1] ^ data_in[7] ^ data_in[6] ^ data_in[1];
    crc_out[7] = crc_reg[15] ^ crc_reg[6] ^ crc_reg[5] ^ crc_reg[0] ^ data_in[6] ^ data_in[5] ^ data_in[0];
    crc_out[6] = crc_reg[14] ^ crc_reg[5] ^ crc_reg[4] ^ data_in[5] ^ data_in[4];
    crc_out[5] = crc_reg[13] ^ crc_reg[7] ^ crc_reg[4] ^ crc_reg[3] ^ crc_reg[1] ^ data_in[7] ^ data_in[4] ^ data_in[3] ^ data_in[1];
    crc_out[4] = crc_reg[12] ^ crc_reg[6] ^ crc_reg[3] ^ crc_reg[2] ^ crc_reg[0] ^ data_in[6] ^ data_in[3] ^ data_in[2] ^ data_in[0];
    crc_out[3] = crc_reg[11] ^ crc_reg[5] ^ crc_reg[2] ^ crc_reg[1] ^ data_in[5] ^ data_in[2] ^ data_in[1];
    crc_out[2] = crc_reg[10] ^ crc_reg[4] ^ crc_reg[1] ^ crc_reg[0] ^ data_in[4] ^ data_in[1] ^ data_in[0];
    crc_out[1] = crc_reg[9] ^ crc_reg[3] ^ crc_reg[0] ^ data_in[3] ^ data_in[0];
    crc_out[0] = crc_reg[8] ^ crc_reg[2] ^ data_in[2];

    return crc_out;
endfunction

function logic [31:0] pre_calc_crc(input logic [7:0] data [0:59]);
    logic [31:0] crc_reg;
    logic [31:0] crc_out;
    integer i;

    crc_reg = 32'hFFFFFFFF;
    for (i = 0; i < 60; i = i + 1) begin
        crc_reg = compute_crc_1(crc_reg, data[i]);
    end

    crc_out = ~crc_reg;

    return crc_out;


endfunction